// memory for computer

module memory(CLK, reset, MemRead, MemWrite, ADDR, Data_in, Data_out);

    reg [15:0] mem[16];
    always@(*) begin
        if (reset)

endmodule